/*
 * generate control signals for 65C02 core.
 *
 * (C) Arlet Ottens <arlet@c-scape.nl>
 */

module ctl(
    input clk,
    input irq,
    input rdy,
    input nmi,
    input reset,
    output sync,
    input cond,
    input [7:0] DB,
    output reg WE,
    output [9:0] flag_op,
    output reg [8:0] alu_op,
    output reg [6:0] reg_op,
    output reg [1:0] do_op,
    output ld_m,
    input I,
    input D,
    output B,
    output reg [11:0] ab_op );

wire [31:0] control;

/*
 * The NMI signal is edge sensitive. Detect edge,
 * register it in 'take_nmi', and clear it at 
 * the next sync pulse, when the NMI is actually
 * taken.
 */
reg nmi1;
reg take_nmi;

always @(posedge clk)
    nmi1 <= nmi;

always @(posedge clk)
    if( nmi & ~nmi1 )
        take_nmi <= 1;
    else if( sync & rdy )
        take_nmi <= 0;

/*
 * take irq when 'irq' is present and not disabled.
 * (priority of irq/nmi will be decided in 'sel_pc' mux)
 */
wire take_irq = irq & ~I;

//assign B = control[8];

reg [3:0] mode;

/*
 * The 4 'mode' bits control the AB datapath. The AB datapath (ABL+ABH) 
 * require a total of 12 control signals, but there are only 15 unique
 * and useful combinations, listed in the table below.
 *
 * The "PC" (consisting of PCH and PCL) is not really the "Program Counter"
 * but simply a holding register for when AB needs to access data. It can
 * either keep the old value, or load it with AB, optionally incremented.
 *
 * The "AHL" is the hold register that stores DB for the next cycle, to be
 * used whenever a 16 bit address appears on the bus. 
 *
 * In case of a branch (mode 0111), the ABL module chooses between DB/00 
 * offset based on its own condition code inputs. The choice for FF/00 
 * for ABH is done here.
 *
 * mode |   PC   | AHL  | AB
 * -----+--------+------+------
 * 0000 |  keep  |  DB  | keep
 * 0001 |  keep  | keep | PC
 * 0010 | AB + 1 |  DB  | {DB, AHL + XYZ} 
 * 0011 | AB + 1 |  DB  | {00, DB  + XYZ} 
 * 0100 |   AB   |  DB  | AB + 1 
 * 0101 |   AB   |  DB  | {01, SP + 1}
 * 0111 |   AB   |  DB  | AB + { FF, DB } + 1   (if backward branch taken) 
 * 0111 |   AB   |  DB  | AB + { 00, DB } + 1   (if forward branch taken)
 * 0111 |   AB   |  DB  | AB + { 00, 00 } + 1   (if branch not taken)
 * 1000 |  keep  | keep | {01, SP} 
 * 1001 | AB + 1 |  DB  | {01, SP}
 * 1010 |  keep  |  DB  | {DB, AHL + XYZ}
 * 1011 |   AB   | keep | {01, SP}
 * 1100 |  keep  |  DB  | AB + 1
 * 1110 |  keep  |  DB  | {DB, AHL + XYZ} + 1
 * 1111 |  keep  | keep | { FF, VECTOR } + 1
 *  |||
 *  |++----> mode bits [1:0] go directly into ABL mux selection
 *  |
 *  +------> mode bit [2] goes directly into ABL carry input
 */

wire abl_ci = mode[2];
wire [1:0] abl_sel = mode[1:0];
wire back = cond & DB[7];     // doing backwards branch 

always @(*)
    case( mode )              //             IPH_ABH____________ABL OP
        4'b0000:                ab_op = { 7'b001_0110, abl_sel, 2'b11, abl_ci };  // AB + 0
        4'b0001:                ab_op = { 7'b000_1010, abl_sel, 2'b10, abl_ci };  // PC
        4'b0010:                ab_op = { 7'b111_1110, abl_sel, 2'b01, abl_ci };  // {DB, AHL+REG}, store PC
        4'b0011:                ab_op = { 7'b111_0000, abl_sel, 2'b01, abl_ci };  // {00, DB+REG}
        4'b0100:                ab_op = { 7'b011_0110, abl_sel, 2'b11, abl_ci };  // AB + 1, store PC
        4'b0101:                ab_op = { 7'b011_0001, abl_sel, 2'b00, abl_ci };  // {01, SP+1}
        4'b0111: if( back )     ab_op = { 7'b011_0111, abl_sel, 2'b11, abl_ci };  // {AB-1, AB} + DB + 1
                 else           ab_op = { 7'b011_0110, abl_sel, 2'b11, abl_ci };  // AB + 1
        4'b1000:                ab_op = { 7'b000_0001, abl_sel, 2'b00, abl_ci };  // {01, SP}, keep PC
        4'b1001:                ab_op = { 7'b111_0001, abl_sel, 2'b00, abl_ci };  // {01, SP}, store PC+1
        4'b1010:                ab_op = { 7'b001_1110, abl_sel, 2'b01, abl_ci };  // {DB, AHL+REG}, keep PC
        4'b1011:                ab_op = { 7'b010_0001, abl_sel, 2'b00, abl_ci };  // {01, SP}
        4'b1100:                ab_op = { 7'b001_0110, abl_sel, 2'b11, abl_ci };  // AB+1, keep PC
        4'b1110:                ab_op = { 7'b001_1110, abl_sel, 2'b01, abl_ci };  // {DB, AHL+REG} + 1, keep PC
        4'b1111:                ab_op = { 7'b000_0011, abl_sel, 2'b00, abl_ci };  // {FF, REG} + 1
        default:                ab_op = { 7'bxxx_xxxx, abl_sel, 2'bxx, abl_ci };  // avoid latches
    endcase

/*
 * control state machine
 */
parameter
    INIT  = 6'd0,
    SYNC  = 6'd1,
    IMM0  = 6'd2,
    IND0  = 6'd3,
    IND1  = 6'd4,
    IND2  = 6'd5,
    DATA  = 6'd6,
    ABS0  = 6'd7,
    ABS1  = 6'd8,
    ZERO  = 6'd9,
    PULL  = 6'd10,
    RDWR  = 6'd11,
    RTS0  = 6'd12,
    RTS1  = 6'd13,
    RTS2  = 6'd14,
    PUSH  = 6'd15,
    JSR0  = 6'd16,
    JSR1  = 6'd17,
    JSR2  = 6'd18,
    BRK0  = 6'd19,
    BRK1  = 6'd20,
    BRK2  = 6'd21,
    BRK3  = 6'd22,
    RTI0  = 6'd23,
    RTI1  = 6'd24,
    RTI2  = 6'd25,
    RTI3  = 6'd26,
    COND  = 6'd27;

reg [5:0] state = INIT;

assign sync = (state == SYNC);

/* 
 * loose state flops
 */
reg rmw, jmp, ind, add_x, add_y, ld, st;
reg [1:0] dst;
reg [3:0] src;
reg [6:0] alu;

/*
 * write enable 
 */
always @(posedge clk)
    case( state )
        BRK0:    WE <= 1;
        BRK1:    WE <= 1;
        BRK2:    WE <= 1;
        JSR0:    WE <= 1;
        JSR1:    WE <= 1;
        PUSH:    WE <= 1;
        RDWR:    WE <= 1;
        default: WE <= 0;
    endcase

/*
 * data output select
 * 
 * 00 ALU
 * 01 P
 * 10 PCL
 * 11 PCH
 */
always @(*)
    case( state )
        BRK1:   do_op = 2'b11;
        BRK2:   do_op = 2'b10;
        BRK3:   do_op = 2'b01;
        JSR1:   do_op = 2'b11;
        JSR2:   do_op = 2'b10;
        DATA:   do_op = 2'b00; 
     default:   do_op = 2'bxx;
    endcase

/*
 * register operation
 *
 *   6   5   4   3   2   1   0
 * +---+---+---+---+---+---+---+
 * | W |  dst  |      src      |
 * +---+---+---+---+---+---+---+
 */
always @(*)
    case( state )
        BRK0:                  reg_op = 7'b1_11_0011; // S
        BRK1:                  reg_op = 7'b1_11_0011; // S
        BRK2:                  reg_op = 7'b1_11_0011; // S
        BRK3:                  reg_op = 7'b0_00_1010; // BRK vector
        JSR0:                  reg_op = 7'b1_11_0011; // S
        JSR1:                  reg_op = 7'b1_11_0011; // S
        RTS0:                  reg_op = 7'b1_11_0011; // S
        RTS1:                  reg_op = 7'b1_11_0011; // S
        RTI0:                  reg_op = 7'b1_11_0011; // S
        RTI1:                  reg_op = 7'b1_11_0011; // S
        RTI2:                  reg_op = 7'b1_11_0011; // S
        PUSH:                  reg_op = 7'b1_11_0011; // S
        PULL:                  reg_op = 7'b1_11_0011; // S
        IND0: if( add_x )      reg_op = 7'b0_00_0000; // X
              else             reg_op = 7'b0_00_0111; // Z
        IND2: if( add_y )      reg_op = 7'b0_00_0001; // Y
              else             reg_op = 7'b0_00_0111; // Z
        ZERO: if( add_x )      reg_op = 7'b0_00_0000; // X
              else if( add_y ) reg_op = 7'b0_00_0001; // Y
              else             reg_op = 7'b0_00_0111; // Z
        ABS1: if( add_x )      reg_op = 7'b0_00_0000; // X
              else if( add_y ) reg_op = 7'b0_00_0001; // Y
              else             reg_op = 7'b0_00_0111; // Z
        SYNC:                  reg_op = { ld, dst, src }; // dst <= src <op> M
        DATA:                  reg_op = { 1'b0, dst, src }; // store
     default:                  reg_op = 7'b0_00_0111; // Z
    endcase

/*
 * ALU operation
 *
 * shift           add
 * -----         --------
 *  10 left      000 OR 
 *  11 right     001 AND
 *               010 XOR
 * carry         011 ADD
 * -----         100 INC
 *  01 1         101 DEC
 *  10 ROT       110 SUB
 *  11 ADC       111 TRB
 *
 *   8   7   6   5   4   3   2   1   0
 * +---+---+---+---+---+---+---+---+---+
 * |ldm|bcd| shift |    add    | carry |
 * +---+---+---+---+---+---+---+---+---+
 */
always @(*)
    case( state )
        BRK0:             alu_op = 9'b00_00_101_00;  // - 1 
        BRK1:             alu_op = 9'b00_00_101_00;  // - 1 
        BRK2:             alu_op = 9'b00_00_101_00;  // - 1 
        JSR0:             alu_op = 9'b00_00_101_00;  // - 1 
        JSR1:             alu_op = 9'b00_00_101_00;  // - 1 
        PUSH:             alu_op = 9'b00_00_101_00;  // - 1
        RTS0:             alu_op = 9'b00_00_100_01;  // + 1 
        RTS1:             alu_op = 9'b00_00_100_01;  // + 1 
        RTI0:             alu_op = 9'b00_00_100_01;  // + 1
        RTI1:             alu_op = 9'b00_00_100_01;  // + 1
        RTI2:             alu_op = 9'b00_00_100_01;  // + 1
        PULL:             alu_op = 9'b00_00_100_01;  // + 1
        IMM0:             alu_op = 9'b10_00_000_00;  // load M
        RDWR:             alu_op = 9'b10_00_000_00;  // load M
        SYNC:             alu_op = {2'b00, alu };    // perform ALU operation
        DATA:    if( st ) alu_op = 9'b00_00_100_00;  // store to M 
                 else     alu_op = {2'b10, alu };    // load M or RMW
        default:          alu_op = 9'bxx_xx_xxx_xx;   
    endcase

always @(*)
    case( state )
        DATA:   mode = 1;
        INIT:   mode = 0;
        SYNC:   mode = 4;
        ABS0:   mode = 4;
        ABS1:   mode = 2;
        IND0:   mode = 3;
        IND1:   mode = 12;
        IND2:   mode = 10;
        ZERO:   mode = 3;
        IMM0:   mode = 4;
        PULL:   mode = 5;
        PUSH:   mode = 11;
        RDWR:   mode = 0;
        RTS0:   mode = 5;
        RTS1:   mode = 5;
        RTS2:   mode = 14;
        RTI0:   mode = 5;
        RTI1:   mode = 5;
        RTI2:   mode = 5;
        RTI3:   mode = 2;
        JSR0:   mode = 9;
        JSR1:   mode = 8;
        JSR2:   mode = 1;
        BRK0:   mode = 9;
        BRK1:   mode = 8;
        BRK2:   mode = 8;
        BRK3:   mode = 15;
        COND:   mode = 7;
    endcase


/*
 * read-modify-write bit. When set, it means
 * we hold the address for extra cycle
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'h06:  rmw <= 1;
            8'hE6:  rmw <= 1;
            8'hEE:  rmw <= 1;
        default:    rmw <= 0;
        endcase

/*
 * jmp bit, indicates that we're jumping to
 * absolute address instead of using it for
 * data
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'h00:  jmp <= 1;
            8'h20:  jmp <= 1;
            8'h40:  jmp <= 1;
            8'h4c:  jmp <= 1;
            8'h60:  jmp <= 1;
            8'h6c:  jmp <= 1;
            8'h7c:  jmp <= 1;
        default:    jmp <= 0;
        endcase

/*
 * indirect bit. Does 16 bit indirected
 * addresses. Needs to be cleared when 
 * used in ABS1 state, otherwise, it will
 * continue to loop indirections.
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'h6c:  ind <= 1;
            8'h7c:  ind <= 1;
        default:    ind <= 0;
        endcase
    else if( state == ABS1 )
        ind <= 0;

/*
 * add_y: use Y register as offset
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'hB1:  add_y <= 1;             // LDA (ZP),Y
            8'hB6:  add_y <= 1;             // LDX ZP,Y
            8'hB9:  add_y <= 1;             // LDX ABS,Y
        default:    add_y <= 0;
        endcase
/*
 * add_x: use X register as offset
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'h7C:  add_x <= 1;             // JMP (IND,X)
            8'hB5:  add_x <= 1;             // LDA ZP,X
            8'hBD:  add_x <= 1;             // LDA ABS,X
            8'hA1:  add_x <= 1;             // LDA (ZP,X)
        default:    add_x <= 0;
        endcase
    else if( state == ABS1 )                // for JMP (IND,X)
        add_x <= 0;

/*
 * ld: load a register at the end of instruction
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'hB1:  ld <= 1;                // LDA (ZP),Y
            8'hB2:  ld <= 1;                // LDA (ZP)
            8'hA1:  ld <= 1;                // LDA (ZP,X)
            8'hA5:  ld <= 1;                // LDA ZP
            8'hA9:  ld <= 1;                // LDA #IMM
            8'hB5:  ld <= 1;                // LDA ZP,X
            8'hAD:  ld <= 1;                // LDA ABS 
            8'hBD:  ld <= 1;                // LDA ABS,X
            8'hB9:  ld <= 1;                // LDA ABS,Y
            8'hB6:  ld <= 1;                // LDX ZP,Y
            8'hA0:  ld <= 1;                // LDY #IMM
            8'hA2:  ld <= 1;                // LDX #IMM
            8'hCA:  ld <= 1;                // DEX 
            8'hE8:  ld <= 1;                // INX
            8'h68:  ld <= 1;                // PLA
        endcase

/*
 * st: store to memory
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'h48:  st <= 1;                // PHA
          default:  st <= 0;        
        endcase

/*
 * src: select source register 
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'hB1:  src <= 7;               // LDA (ZP),Y
            8'hB2:  src <= 7;               // LDA (ZP)
            8'hA1:  src <= 7;               // LDA (ZP,X)
            8'hA5:  src <= 7;               // LDA ZP
            8'hA9:  src <= 7;               // LDA #IMM
            8'hB5:  src <= 7;               // LDA ZP,X
            8'hAD:  src <= 7;               // LDA ABS 
            8'hBD:  src <= 7;               // LDA ABS,X
            8'hB9:  src <= 7;               // LDA ABS,Y
            8'hA2:  src <= 7;               // LDX #IMM 
            8'hB6:  src <= 7;               // LDX ZP,Y
            8'hCA:  src <= 0;               // DEX 
            8'hE8:  src <= 0;               // INX
            8'h68:  src <= 7;               // PLA
            8'h48:  src <= 2;               // PHA 
            8'hA0:  src <= 7;               // LDY #IMM 
            8'hE6:  src <= 5;               // INC ZP
            8'hEE:  src <= 5;               // INC ABS 
        endcase

/*
 * dst: select destination register 
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'hB1:  dst <= 2;               // LDA (ZP),Y
            8'hB2:  dst <= 2;               // LDA (ZP)
            8'hA1:  dst <= 2;               // LDA (ZP,X)
            8'hA5:  dst <= 2;               // LDA ZP
            8'hA9:  dst <= 2;               // LDA #IMM
            8'hB5:  dst <= 2;               // LDA ZP,X
            8'hAD:  dst <= 2;               // LDA ABS 
            8'hBD:  dst <= 2;               // LDA ABS,X
            8'hB9:  dst <= 2;               // LDA ABS,Y
            8'h68:  dst <= 2;               // PLA

            8'hA2:  dst <= 0;               // LDX #IMM 
            8'hB6:  dst <= 0;               // LDX ZP,Y
            8'hCA:  dst <= 0;               // DEX 
            8'hE8:  dst <= 0;               // INX

            8'hA0:  dst <= 1;               // LDY #IMM 
        endcase

/*
 * alu: select ALU operation 
 */
always @(posedge clk)
    if( sync )
        case( DB )
            8'hB1:  alu <= 7'b00_011_00;    // LDA (ZP),Y
            8'hB2:  alu <= 7'b00_011_00;    // LDA (ZP)
            8'hA1:  alu <= 7'b00_011_00;    // LDA (ZP,X)
            8'hA5:  alu <= 7'b00_011_00;    // LDA ZP
            8'hA9:  alu <= 7'b00_011_00;    // LDA #IMM
            8'hB5:  alu <= 7'b00_011_00;    // LDA ZP,X
            8'hAD:  alu <= 7'b00_011_00;    // LDA ABS 
            8'hBD:  alu <= 7'b00_011_00;    // LDA ABS,X
            8'hB9:  alu <= 7'b00_011_00;    // LDA ABS,Y
            8'hA2:  alu <= 7'b00_011_00;    // LDX #IMM 
            8'hB6:  alu <= 7'b00_011_00;    // LDX ZP,Y
            8'hA0:  alu <= 7'b00_011_00;    // LDY #IMM 

            8'hCA:  alu <= 7'b00_101_00;    // DEX 
            8'hE8:  alu <= 7'b00_100_01;    // INX

            8'hE6:  alu <= 7'b00_011_00;    // INC ZP
            8'hEE:  alu <= 7'b00_011_00;    // INC ABS 
            
            8'h48:  alu <= 7'b00_011_00;    // PHA
            8'h68:  alu <= 7'b00_011_00;    // PLA
        default:    alu <= 7'b11_111_11;    // don't care
        endcase

always @(posedge clk)
    case( state )
        INIT:   state <= SYNC;
        SYNC:   
            case( DB )
                8'h80:  state <= COND;      // BRA
                8'h00:  state <= BRK0;      // BRK
                8'h20:  state <= JSR0;      // JSR
                8'h40:  state <= RTI0;      // RTI
                8'h60:  state <= RTS0;      // RTS
                8'h4C:  state <= ABS0;      // JMP ABS
                8'h6C:  state <= ABS0;      // JMP (IND)
                8'h7C:  state <= ABS0;      // JMP (IND,X)
                8'h06:  state <= ZERO;      // ASL ZP
                8'h16:  state <= ZERO;      // ASL ZP,X
                8'hA5:  state <= ZERO;      // LDA ZP
                8'hB5:  state <= ZERO;      // LDA ZP,X
                8'hB6:  state <= ZERO;      // LDX ZP,Y
                8'hA1:  state <= IND0;      // LDA (ZP,X)
                8'hB2:  state <= IND0;      // LDA (ZP)
                8'hB1:  state <= IND0;      // LDA (ZP),Y
                8'hAD:  state <= ABS0;      // LDA ABS 
                8'hBD:  state <= ABS0;      // LDA ABS,X
                8'hB9:  state <= ABS0;      // LDA ABS,Y
                8'hA9:  state <= IMM0;      // LDA #IMM
                8'hA0:  state <= IMM0;      // LDY #IMM
                8'hA2:  state <= IMM0;      // LDX #IMM
                8'h48:  state <= PUSH;      // PUSH
                8'h68:  state <= PULL;      // PULL
                8'hE6:  state <= ZERO;      // INC ZP
                8'hEE:  state <= ABS0;      // INC ABS 
            endcase
        IND0:   state <= IND1;
        IND1:   state <= IND2;      //
        IND2:   state <= DATA;
        IMM0:   state <= SYNC;
        ABS0:   state <= ABS1;
        ZERO:   state <= rmw ? RDWR : DATA;
        ABS1:   state <= ind ? ABS0 : 
                         jmp ? SYNC : 
                         rmw ? RDWR : DATA;
        RDWR:   state <= DATA;
        DATA:   state <= SYNC;
        PULL:   state <= DATA;
        PUSH:   state <= DATA;
        RTS0:   state <= RTS1;
        RTS1:   state <= RTS2;
        RTS2:   state <= SYNC; 
        JSR0:   state <= JSR1;
        JSR1:   state <= JSR2;
        JSR2:   state <= ABS1;
        BRK0:   state <= BRK1;
        BRK1:   state <= BRK2;
        BRK2:   state <= BRK3;
        BRK3:   state <= ABS0;
        RTI0:   state <= RTI1;
        RTI1:   state <= RTI2;
        RTI2:   state <= RTI3;
        RTI3:   state <= SYNC;
        COND:   state <= SYNC;
    endcase

`ifdef SIM
reg [31:0] statename;

always @(*)
    case( state )
        INIT: statename = "INIT";
        SYNC: statename = "SYNC";
        DATA: statename = "DATA";
        IMM0: statename = "IMM0";
        DATA: statename = "DATA";
        IND0: statename = "IND0";
        IND1: statename = "IND1";
        IND2: statename = "IND2";
        ABS0: statename = "ABS0";
        ABS1: statename = "ABS1";
        PULL: statename = "PULL";
        PUSH: statename = "PUSH";
        ZERO: statename = "ZERO";
        RDWR: statename = "RDWR";
        RTS0: statename = "RTS0";
        RTS1: statename = "RTS1";
        RTS2: statename = "RTS2";
        JSR0: statename = "JSR0";
        JSR1: statename = "JSR1";
        JSR2: statename = "JSR2";
        BRK0: statename = "BRK0";
        BRK1: statename = "BRK1";
        BRK2: statename = "BRK2";
        BRK3: statename = "BRK3";
        RTI0: statename = "RTI0";
        RTI1: statename = "RTI1";
        RTI2: statename = "RTI2";
        RTI0: statename = "RTI3";
        COND: statename = "COND";
    endcase
`endif

endmodule
